`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/08/2021 04:25:18 PM
// Design Name: 
// Module Name: LinearInterpolator
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
//
// Additional Comments:
//  Interpolation formular: InterpValue = snd_data[1]*(maxCnt - smplCnt) + snd_data[0]*(smplCnt)
//                          InterpValue = snd_data[1]*(sub_sample_count - intrp_sub_sample) + snd_data[0]*intrp_sub_sample
//
//
//                           InterpValue
//                               V
//                      X--------|--------------X               >> time, X = input sample points
//               snd_data[1]                snd_data[0]         >> V = 96KHz sample points
//                      |<--a--->|
//                      |<------- maxCnt -------|
//////////////////////////////////////////////////////////////////////////////////
//
//      


module LinearInterpolator(
    input           clk,
    input           reset_n,
    input           run,
    input           l_din_en,      // ignore and just use r_din_en for both channels
    input           r_din_en,
    input [23:0]    l_data_in,
    input [23:0]    r_data_in,
 //   input [9:0]     sub_sample_cnt,
    output reg      dout_valid,
    output [33:0]   l_data_out,
    output [33:0]   r_data_out,
    // for test
    output reg [2:0]   interp_state,
    input [1:0]     test_d_select,
    output [15:0]    test_data 
);

reg [1:0]   l_snd_data[23:0];
reg [1:0]   r_snd_data[23:0];
reg [1:0]   l_intrp_data[23:0];
reg [1:0]   r_intrp_data[23:0];
reg [1:0]   intrp_coef[9:0];
reg [9:0]   mult_coef;
reg         mult_en, dout_en, coef_sub_en, adder_en;
// reg [2:0]   interp_cnt;
reg [23:0]  l_mult_din, r_mult_din;
reg [33:0]  l_mult_dout, r_mult_dout;
reg [1:0]   l_dout[32:0];
reg [1:0]   r_dout[32:0];
reg [9:0]   input_max_sample_count, input_sample_count, input_sample_counter; 
reg [9:0]   intrp_input_count, intrp_input_max_count;
reg [10:0]  sample_1_coef, sample_96KHz_count;


parameter sample_96KHz_max = 10'h1ff;      // divide by 512 for 96KHz (programmabe later?)



// generate System sample clk @ 96KHz
// divide mclk 49.152MHz by sample_96KHz_max (512) to create 96000Hz
always @ (posedge clk) begin
    if (!run) begin
        dout_en <= 1'b0;
        sample_96KHz_count <= 0;
        input_sample_count <= 0;
    end
    else if (sample_96KHz_count == sample_96KHz_max) begin
        sample_96KHz_count <= 0;
        dout_en <= 1'b1;
        input_sample_count <= input_sample_counter;     // hold count value at the 96KHz sample
    end
    else begin
        sample_96KHz_count <= sample_96KHz_count + 1;
        dout_en <= 1'b0;
        input_sample_count <= input_sample_count;
    end
end

// Capture Input Data
// access 2 consecutive samples (l & r) and sub_sample count between the 2 samples
// get coefficient from sub sample count
always @ (posedge clk) begin
    if(r_din_en) begin              // strobe, start/end of a sample
        input_sample_counter <= 0;
        r_snd_data[0] <= r_data_in;
        r_snd_data[1] <= r_snd_data[0];
        l_snd_data[0] <= l_data_in;
        l_snd_data[1] <= l_snd_data[0];
        input_max_sample_count <= input_sample_counter;
    end
    else begin
        input_sample_counter <= input_sample_counter + 1;        
        r_snd_data <= r_snd_data;
        l_snd_data <= l_snd_data;
        input_max_sample_count <= input_max_sample_count; 
    end
end           

// Hold Input Data if State Machine Active
always @ (posedge clk) begin
    if(interp_state == 0) begin               
        l_intrp_data <= l_snd_data;
        r_intrp_data <= r_snd_data;
        intrp_input_count <= input_sample_count;            // 96KHz position relative to input sample  (a)
        intrp_input_max_count <= input_max_sample_count;    // total mclks between input samples        (1)
    end
    else begin
        l_intrp_data <= l_intrp_data;
        r_intrp_data <= r_intrp_data;
        intrp_input_count <= intrp_input_count;
        intrp_input_max_count <= intrp_input_max_count;
    end
end

    

// Interpolatator State Machine
always @ (posedge clk) begin
    case (interp_state)
        0: begin
            mult_en <= 1'b0;
            dout_valid <= 1'b0;
            intrp_coef <= intrp_coef;
            
            if (dout_en) begin  
                interp_state <= 1;
                coef_sub_en <= 1;       // enable subtractor
            end
            else begin
                interp_state <= 0;
                coef_sub_en <= 0;
            end
        end
        1: begin
            interp_state <= 2;
            mult_en <= 1'b0;
            dout_valid <= 1'b0;
            // prevent a negative number
            if (sample_1_coef[10]) begin // if the result is negative, then a = intrp_input_max_count
                intrp_coef[1] <= 0;                         // a-a=0
                intrp_coef[0] <= intrp_input_max_count;     // a=1
            end
            else begin
                intrp_coef[1] <= sample_1_coef[9:0];        // subtracter result:  1 - a 
                intrp_coef[0] <= intrp_input_count;         // max input samples:  a
            end
        end
            
        2: begin
            interp_state <= 3;
            mult_en <= 1'b0;
            dout_valid <= 1'b0;
            l_mult_din <= l_intrp_data[0];
            r_mult_din <= r_intrp_data[0];
            mult_coef <= intrp_coef[0];
        end
        
        3: begin
            interp_state <= 4;
            mult_en <= 1'b1;
            dout_valid <= 1'b0;
            l_mult_din <= l_intrp_data[1];
            r_mult_din <= r_intrp_data[1];
            mult_coef <= intrp_coef[1];
           
        end    
        4: begin
            interp_state <= 5;
            mult_en <= 1'b1;
            dout_valid <= 1'b0;
            l_dout[0] <= l_mult_dout[33:1];
            r_dout[0] <= r_mult_dout[33:1];
        end
        5: begin
            interp_state <= 6;
            mult_en <= 1'b0;
            adder_en <= 1'b1;
            dout_valid <= 1'b0;
            l_dout[1] <= l_mult_dout[33:1];
            r_dout[1] <= r_mult_dout[33:1];
        end         
        6: begin
            interp_state <= 0;
            mult_en <= 1'b0;
            adder_en <= 1'b0;
            dout_valid <= 1'b1;            
        end
        default: begin
            mult_en <= 1'b0;
            adder_en <= 1'b0;
            dout_valid <= 1'b0;
            interp_state <= 0;
            intrp_coef <= intrp_coef;
        end
    endcase
end
                

interpolator_subtractor l_interp_sub (
    .A            (intrp_input_max_count),  // input wire [9 : 0] A
    .B            (intrp_input_count),      // input wire [9 : 0] B
    .CLK          (clk),                    // input wire CLK
    .CE           (coef_sub_en),            // input wire CE
    .S            (sample_1_coef)           // output wire [10 : 0] S
);

                

interp_mult l_interp_mult (
    .CLK    (clk),              // input wire CLK
    .CE     (mult_en),          // input wire CE
    .A      (l_mult_din),       // input wire [23 : 0] B
    .B      (mult_coef),        // input wire [9 : 0] A
    .P      (l_mult_dout)       // output wire [33 : 0] P);
 );
   
interp_mult r_interp_mult (
    .CLK    (clk),              // input wire CLK
    .CE     (mult_en),          // input wire CE
    .A      (r_mult_din),       // input wire [23 : 0] B
    .B      (mult_coef),        // input wire [9 : 0] A
    .P      (r_mult_dout)       // output wire [33 : 0] P);
 );
   
Interpolator_adder l_interp_add (
  .A            (l_dout[0]),            // input wire [32 : 0] A
  .B            (l_dout[1]),            // input wire [32 : 0] B
  .CLK          (clk),                  // input wire CLK
  .CE           (add_en),               // input wire CE
  .S            (l_data_out)            // output wire [33 : 0] S
);

Interpolator_adder r_interp_add (
  .A            (r_dout[0]),            // input wire [32 : 0] A
  .B            (r_dout[1]),            // input wire [32 : 0] B
  .CLK          (clk),                  // input wire CLK
  .CE           (add_en),               // input wire CE
  .S            (r_data_out)            // output wire [33 : 0] S
);


//      TEST


assign test_data =      (test_d_select == 0) ?  r_data_in[15:0] :
                        (test_d_select == 1) ?  r_data_in[23:8] :
                        (test_d_select == 2) ?  l_data_in[15:0] :
                                                l_data_in[23:8];

endmodule
